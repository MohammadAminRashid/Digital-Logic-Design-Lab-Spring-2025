module const8bit(
    output [7:0] val
);
    assign val = 8'b00000000;
endmodule